module accelerator #(
    globalBufferSize = 1024,
    globalBufferInterfaceSize = 16,
    dataSize = 8
) (
    
);
    
// Global Buffer Interface


endmodule