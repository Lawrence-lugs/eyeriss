module accelerator #(
    globalBufferSize = 1024,
    dataSize = 8,
    globalBufferInterfaceSize =  
) (
    
);
    
// Global Buffer Interface


endmodule